// ula_opcodes.vh
`define ADD   4'b0000
`define SUB   4'b0001
`define AND   4'b0010
`define OR    4'b0011
`define XOR   4'b0100
`define NOR   4'b0101
`define SLT   4'b0110
`define SLTU  4'b0111
`define SLL   4'b1000
`define SRL   4'b1001
`define SRA   4'b1010
`define SLLV  4'b1011
`define SRLV  4'b1100
`define SRAV  4'b1101
`define JR    4'b1110
